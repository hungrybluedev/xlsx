module xlsx

// pub fn (sheet Sheet) get_cell

module xlsx

// Sets a string cell at the given location
pub fn (mut sheet Sheet) set_cell(loc Location, value string) {
	sheet.ensure_row_exists(loc.row)
	row_idx := sheet.find_row_index(loc.row)
	sheet.rows[row_idx].cells << Cell{
		cell_type: .string_type
		location:  loc
		value:     value
	}
}

// Sets a numeric cell at the given location (int version)
pub fn (mut sheet Sheet) set_number(loc Location, value int) {
	sheet.ensure_row_exists(loc.row)
	row_idx := sheet.find_row_index(loc.row)
	sheet.rows[row_idx].cells << Cell{
		cell_type: .number_type
		location:  loc
		value:     value.str()
	}
}

// Sets a numeric cell at the given location (f64 version)
pub fn (mut sheet Sheet) set_number_f64(loc Location, value f64) {
	sheet.ensure_row_exists(loc.row)
	row_idx := sheet.find_row_index(loc.row)
	sheet.rows[row_idx].cells << Cell{
		cell_type: .number_type
		location:  loc
		value:     value.str()
	}
}

// Sets a formula cell at the given location
pub fn (mut sheet Sheet) set_formula(loc Location, formula string) {
	sheet.ensure_row_exists(loc.row)
	row_idx := sheet.find_row_index(loc.row)
	sheet.rows[row_idx].cells << Cell{
		cell_type: .number_type // Formulas are typically numbers
		location:  loc
		value:     '' // Value will be computed by Excel
		formula:   formula
	}
}

// Ensures a row exists at the given index, creating it if necessary
fn (mut sheet Sheet) ensure_row_exists(row_index int) {
	// Check if row already exists
	for r in sheet.rows {
		if r.row_index == row_index {
			return
		}
	}
	// Create new row
	sheet.rows << Row{
		row_index: row_index
		row_label: (row_index + 1).str()
		cells:     []Cell{}
	}
}

// Finds the internal index of a row by its row_index
fn (sheet Sheet) find_row_index(row_index int) int {
	for i, r in sheet.rows {
		if r.row_index == row_index {
			return i
		}
	}
	return -1 // Should not happen if ensure_row_exists was called
}
